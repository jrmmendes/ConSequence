-------------------------------------------------
-- Contador parametrizado
-- Por Jose R. M. Junior <jrmmendes@outlook.com>
-- Ultima modificacao: 09/10/2018 11:52
-------------------------------------------------
-- Bibliotecas ----------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Entidade -------------------------------------
entity NomeDaEntidade is
  generic(
  -- parametros
  );
  port(
  -- portas
  );
end entity;
-- Arquiteturas ---------------------------------
architecture nomeDaArquitetura of NomeDaEntidade is

begin
  -- descricao comportamental
end architecture;